// list all paths to your design files
`include "../PE_array_64.v"
`include "../PE.v"
`include "../memory_control.v"